PACKAGE Common IS
	TYPE state_type IS (idle, loadRNG, enableRNG, loadSR, transmit);
END Common;